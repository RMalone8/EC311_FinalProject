`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/08/2023 02:31:20 PM
// Design Name: 
// Module Name: WordLibrary
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module WordDelivery(
    clk,
    wordComplete,
    reset,
    
    currentWord,
    nextWord
    );
    
input clk;
input wordComplete;
input reset;

output reg [19:0] currentWord;
output reg [19:0] nextWord;
 
reg [19:0] word [0:99];
wire [6:0] nextWordLocation;

RandomNumberGenerator randomizer(.grabWord(wordComplete), .reset(reset), .random_num(nextWordLocation));

always @ (posedge wordComplete) begin
    currentWord = nextWord;
    nextWord = word[nextWordLocation];
end




initial begin
    
    word[0] = 20'b00001100100000010111;
    word[1] = 20'b00010101010000000001;
    word[2] = 20'b01010100100101100100;
    word[3] = 20'b01111100101001001011;
    word[4] = 20'b00010000000111101111;
    word[5] = 20'b00011100100011110110;
    word[6] = 20'b10011100101010101011;
    word[7] = 20'b10101100101001010000;
    word[8] = 20'b10111001000001001000;
    word[9] = 20'b00000011111011010010;
    word[10] = 20'b11101001001011010111;
    word[11] = 20'b11100000001010110001;
    word[12] = 20'b10100110000100110011;
    word[13] = 20'b01010010011000111011;
    word[14] = 20'b11010001000111100011;
    word[15] = 20'b10010001110111100100;
    word[16] = 20'b10000001000111100011;
    word[17] = 20'b01111110001011001000;
    word[18] = 20'b01011010011011100100;
    word[19] = 20'b01010100100111110111;
    word[20] = 20'b01000000001110111100;
    word[21] = 20'b00111110001011001000;
    word[22] = 20'b00101011110000001011;
    word[23] = 20'b00100000100100010010;
    word[24] = 20'b00011110001011001011;
    word[25] = 20'b00010110001011010011;
    word[26] = 20'b00001011110100110011;
    word[27] = 20'b00000110001010100000;
    word[28] = 20'b00000100110010011011;
    word[29] = 20'b11010010011011010011;
    word[30] = 20'b11001001000100101111;
    word[31] = 20'b11000100010001110010;
    word[32] = 20'b10111000000001010111;
    word[33] = 20'b10110110100100100111;
    word[34] = 20'b10101110000000111100;
    word[35] = 20'b10011010011011101000;
    word[36] = 20'b10010100110000001111;
    word[37] = 20'b10000110001011000100;
    word[38] = 20'b01111100100000100100;
    word[39] = 20'b01011010011101001001;
    word[40] = 20'b01001101010100110110;
    word[41] = 20'b01000000000111110010;
    word[42] = 20'b00111000001110100100;
    word[43] = 20'b00101010011110111101;
    word[44] = 20'b00100100110100100010;
    word[45] = 20'b00011110001000100100;
    word[46] = 20'b00010011110000011010;
    word[47] = 20'b00001101010100110000;
    word[48] = 20'b00000110010100100011;
    word[49] = 20'b11010000001000100100;
    word[50] = 20'b10111101010010001011;
    word[51] = 20'b10110100001100000111;
    word[52] = 20'b10101010010010110111;
    word[53] = 20'b10011011111001000011;
    word[54] = 20'b00000110110111100100;
    word[55] = 20'b00001000000111110000;
    word[56] = 20'b00010010001100000111;
    word[57] = 20'b00011100101000000100;
    word[58] = 20'b00100100011100111100;
    word[59] = 20'b00101000001000100111;
    word[60] = 20'b00111011111100000100;
    word[61] = 20'b01000110001011001000;
    word[62] = 20'b01001000111001001111;
    word[63] = 20'b01010000000001001011;
    word[64] = 20'b01011001000010010001;
    word[65] = 20'b01111010011000010011;
    word[66] = 20'b10000110001011100100;
    word[67] = 20'b10001100101001001011;
    word[68] = 20'b10010000001011101000;
    word[69] = 20'b10011001000000001011;
    word[70] = 20'b10101110001011000100;
    word[71] = 20'b10110010010010110111;
    word[72] = 20'b10111100101010110001;
    word[73] = 20'b11000101010011100100;
    word[74] = 20'b11001000001011010111;
    word[75] = 20'b11010000001010110011;
    word[76] = 20'b11011111001011010111;
    word[77] = 20'b11100001000111110011;
    word[78] = 20'b11101100101000100100;
    word[79] = 20'b00000000010010010111;
    word[80] = 20'b00001100100111110111;
    word[81] = 20'b00010110000111101111;
    word[82] = 20'b00011000001000010011;
    word[83] = 20'b00100000001010101111;
    word[84] = 20'b00101000000001100100;
    word[85] = 20'b00111101010100110111;
    word[86] = 20'b01000001001010100001;
    word[87] = 20'b01001000100010000011;
    word[88] = 20'b01010100101101001111;
    word[89] = 20'b01011100010100110111;
    word[90] = 20'b01111000001010101011;
    word[91] = 20'b10000010011010100100;
    word[92] = 20'b10001000001001100100;
    word[93] = 20'b10010100101110100100;
    word[94] = 20'b10011110000001001011;
    word[95] = 20'b10101100100000010000;
    word[96] = 20'b10110001000010010011;
    word[97] = 20'b10111110001011001011;
    word[98] = 20'b11000011111000100000;
    word[99] = 20'b11001001000010010101;
end

endmodule