`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/08/2023 02:31:20 PM
// Design Name: 
// Module Name: WordLibrary
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module WordDelivery(
    clk,
    wordComplete,
    reset,
    
    currentWord,
    nextWord
    );
    
input clk;
input wordComplete;
input reset;

output reg [19:0] currentWord;
output reg [19:0] nextWord;
 
reg [19:0] word [0:99];
wire [6:0] nextWordLocation;

RandomNumberGenerator randomizer(.grabWord(wordComplete), .reset(reset), .random_num(nextWordLocation));

always @ (posedge wordComplete) begin
    currentWord = nextWord;
    nextWord = word[nextWordLocation];
end




initial begin
    
    word[0] = 20'b00001011100000010011;
    word[1] = 20'b00010100010000000001;
    word[2] = 20'b01001011100101000100;
    word[3] = 20'b01011011100111001010;
    word[4] = 20'b00010000000101101011;
    word[5] = 20'b00011011100011010010;
    word[6] = 20'b01111011101000101010;
    word[7] = 20'b10001011100111001100;
    word[8] = 20'b10011001000001000111;
    word[9] = 20'b00000010111001001110;
    word[10] = 20'b11001001001001010011;
    word[11] = 20'b11000000001000101101;
    word[12] = 20'b10000101000100001111;
    word[13] = 20'b01001010000110110111;
    word[14] = 20'b10110001000101100011;
    word[15] = 20'b01110001100101100100;
    word[16] = 20'b01100001000101100011;
    word[17] = 20'b01011101001001000111;
    word[18] = 20'b01010010001001100100;
    word[19] = 20'b01001011100101110011;
    word[20] = 20'b00111000001100111000;
    word[21] = 20'b00110101001001000111;
    word[22] = 20'b00101010110000001010;
    word[23] = 20'b00100000100011101110;
    word[24] = 20'b00011101001001001010;
    word[25] = 20'b00010101001001001111;
    word[26] = 20'b00001010110100001111;
    word[27] = 20'b00000101001000100000;
    word[28] = 20'b00000011110010010111;
    word[29] = 20'b10110010001001001111;
    word[30] = 20'b10101001000100001011;
    word[31] = 20'b10100011010001101110;
    word[32] = 20'b10011000000001010011;
    word[33] = 20'b10010101100100000110;
    word[34] = 20'b10001101000000111000;
    word[35] = 20'b01111010001001100111;
    word[36] = 20'b01110011110000001011;
    word[37] = 20'b01100101001001000100;
    word[38] = 20'b01011011100000100100;
    word[39] = 20'b01010010001011001000;
    word[40] = 20'b01000100010100010010;
    word[41] = 20'b00111000000101101110;
    word[42] = 20'b00110000001100100100;
    word[43] = 20'b00101010001100111001;
    word[44] = 20'b00100011110100000010;
    word[45] = 20'b00011101000110100100;
    word[46] = 20'b00010010110000010110;
    word[47] = 20'b00001100010100001100;
    word[48] = 20'b00000101010100000011;
    word[49] = 20'b10110000000110100100;
    word[50] = 20'b10011100010010001010;
    word[51] = 20'b10010011001010000110;
    word[52] = 20'b10001010000010110011;
    word[53] = 20'b01111010110111000011;
    word[54] = 20'b00000101110101100100;
    word[55] = 20'b00001000000101101100;
    word[56] = 20'b00010001111010000110;
    word[57] = 20'b00011011100110000100;
    word[58] = 20'b00100011011010111000;
    word[59] = 20'b00101000000110100110;
    word[60] = 20'b00110010111010000100;
    word[61] = 20'b00111101001001000111;
    word[62] = 20'b01000000110111001011;
    word[63] = 20'b01001000000001001010;
    word[64] = 20'b01010001000010001101;
    word[65] = 20'b01011010000110001111;
    word[66] = 20'b01100101001001100100;
    word[67] = 20'b01101011100111001010;
    word[68] = 20'b01110000001001100111;
    word[69] = 20'b01111001000000001010;
    word[70] = 20'b10001101001001000100;
    word[71] = 20'b10010010000010110011;
    word[72] = 20'b10011011101000101101;
    word[73] = 20'b10100100010011000100;
    word[74] = 20'b10101000001001010011;
    word[75] = 20'b10110000001000101111;
    word[76] = 20'b10111110001001010011;
    word[77] = 20'b11000001000101101111;
    word[78] = 20'b11001011100110100100;
    word[79] = 20'b00000000010010010011;
    word[80] = 20'b00001011100101110011;
    word[81] = 20'b00010101000101101011;
    word[82] = 20'b00011000000110001111;
    word[83] = 20'b00100000001000101011;
    word[84] = 20'b00101000000001100100;
    word[85] = 20'b00110100010100010011;
    word[86] = 20'b00111001001000100001;
    word[87] = 20'b01000000100010000011;
    word[88] = 20'b01001011101011001011;
    word[89] = 20'b01010011010100010011;
    word[90] = 20'b01011000001000101010;
    word[91] = 20'b01100010001000100100;
    word[92] = 20'b01101000000111100100;
    word[93] = 20'b01110011101100100100;
    word[94] = 20'b01111101000001001010;
    word[95] = 20'b10001011100000001100;
    word[96] = 20'b10010001000010001111;
    word[97] = 20'b10011101001001001010;
    word[98] = 20'b10100010110110100000;
    word[99] = 20'b10101001000010010001;
end

endmodule